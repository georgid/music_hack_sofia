BZh91AY&SY��*w �_�Py��g߰����P��dqؖl���(�SdS�1G��4��i��4424@�C$�D =M�    ��B��i<��O�C�Ʉ`�h{E4�sbh0�2d��`�i���!�IA4�Ҟ�G��i�2=@  4hRC�! V@���(�߀�}�f�m�(#G�O�f	!�.��hv7p��졪�d\���G��D��:��c(�7�eF���̇g��v���� ɖ��Ю�0�)��G C,t�S}�B��H�@�ʌ�E�,�})��$� �d0׾�n�C�̲G\�-l�\�1���!�B�8���l�c{^��q<��Qr�39�Vƣ仆��z���w�-$D\�Z�$��"Sx��Q&�%��16��*�i�2��Su��EF�Km��С /�.P�3�Ĳ�R���p�{��e�s&%�A_P�P���K@[����R��ճ�Xzu3���H�#c7L���G�h�/H4�M-���-L���� �)V�O�W4����qp��+��[�aC��iQb>�0%*j�[E�f�6�4�=
�`0C�vC{:��@:������v�]�������݃k"�P�i���J��:������ݏZI�־*��o���:�"9���W���x5 �G(�m
�0
�[S�aT��䂤r�Td;�d	�>rz�LRFw��PZ�w��R�ʩ0i��>�-�\g����S��r���淸?����\tb�����	v�^�}�Ê�Q��N�&�l�0nᘨR�QhO�AsF@��Ʃ�|�
��N��=�LŉЀȽ��:X�̋ܒ���I�d���l�a��32�׀>�[�B�aG>;
H��<�A�{X$f,���Й��u��q5'"�'	��R��y�� �=D�=;n-N�ݓ'<A���)A�<0��QC�Ũ��O=u�`@���'�vETP����%��5��=�p�����4��:feD�c�0m�@��B렘��3s���j_-�Qĥ��;��J�D�D,ˁ S�h����\FA��=�VѨ)��l�4	��AYYk��yqR_
+����Co��͢+]���>���s�`�Ԍ��w$S�	
|��p