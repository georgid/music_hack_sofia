BZh91AY&SY�e� �߀Ry����������`	|>����d �� )F���zC  ��  �i%��     �#!�4a0F�4b�20 I���M)��`��4���Pdh�sL��Lф�hшd�� A"D�#�$���<�Mi��i�4z����;0��Ԓ�hd&I!
 ��zF,�k�O8���Y���w�z��g2Dd��5 �=A�´L�H@�%ň~��5?j*������4ha�����O����9�r ��.�VF��!;�u#�sF�I�]����8@�	�a�����TJt�Ғ�d�j�⚪DNQ~g�/��ɶSa/n�1� f�i�,�
	O�)R1�de�VDP��k,1��fY�w��y�,8�)�<�3<u걕�o��I"���"_gc�W�[��
�#p^v���1/.m���2/1�8�KE2���X����CM���9�L�Yލ�TA�#�T�Sņ�z�	�&@Q=e�H�K���a��p��ny�׉���7��`���U����L�d}FR
�	4b��rfɓ�����ݺ]��M)���Uq�tTh�/�Ȳ���d0{��= F���K)7�i.J��],�<.�E��C�ɐ�A������*����@hZjr����0)�R���0��Z*��m��"-E�ұ�����E�AmA�2d�)�g�U��U欘F!��"(a�D���yy�e< C.wiY%0��Ӈ����J�$j�!CVPP���� ��hĘYKC�a���ˉ��	������N���J��$8;=O��DԬ`yX}�J�6�їA��2�z�*��UB�pE�E��k	�;�ɤ-+kK�?9r����fŧ�Ƙ9���%D8��l�PZl����I�ܠ���N5w���@*��rNIɦ����W�����0�n4{�ȩ���Y��.��}���?#�2�AEԁ�7t���������A;����+��d*B���ffZu�tO��ɅĪ��\L�W��N�A�F���l@�?`�|g�������-i
��4h�B!"G���l�xg��6��U� &�s�T��s�\�%�3���7���B�K�B����+�5Z�
�0��z�R|2�6��bU�� ��hH,VNħq9�L�E�lo15���;��H����I���4���}Nc��u/!�\�%܈��J ���1Lb�,+0��m���9�A�� �V�EM�`i]��`"I�QiMx���,UX4��D	�F��-�-(�3�3Jх�t5h���PG}��8��� ���\�@5d�BIoJeR����N{��/�ZJ�qa�%"S�$�E�{��]�ys.%Q���z��yA���d��ܟj,:�]�h��DA�m��z й�1��I� `���s�'w:�B�H�/yy%�/%����_�Ĩ3Rb�K[@�~��3^�5�s^EW'ɱ2`^3��!�UsF�*C���v'�h�\�Ԛ��1�r,J,�AQ7�碈H��YӿD�O�f@�.p�
"FJjI��'l�!�6g �-� ��D�`i��V0���|KRLaq~K��v��}%B�u����U#Ӹ�xl70C���J�.�_1�	�} +�APl��\ ��$))P��Mr�E�>�ؗp��1�8�V���W�y������ 	��6̭Y9�u��C5�	M��%!TrJG�nk� ���X�<ϩ^�j&^z�P��5$��\�
DQ!�$uj%Φ�1��b$�|�-���KS.\��.��8�%AA��5&�-6�I�I@����0��X��Ъ�:	�5kg1Tq�9��)!���-L S�25"ĵ�w^���
�C#J�5�I�(k�̺�L��m�6Դ&�n����w��/��͠i�U<	��=����1��Q#��#�a���Áp`�����8p�tEJ�
��	���+o����od����p J�խ?�]��BC����